module Picture_Shifter (
    input clk,
    input rst,
    input random_num,
    input shift,
    input Gaming,
    input ready,
    output R0in,
    output R1in,
    output B0in,
    output B1in,
    output G0in,
    output G1in,
);
    

    
endmodule

module matrix_generate(
    input clk,
    input rst, 
    input col,
    input row,
    output R0,
    output B0,
    output G0,
    output R1,
    output B1,
    output G1
);

